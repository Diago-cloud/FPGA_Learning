library verilog;
use verilog.vl_types.all;
entity TB_Seq_101 is
end TB_Seq_101;
