library verilog;
use verilog.vl_types.all;
entity TB_LED_PWM is
end TB_LED_PWM;
